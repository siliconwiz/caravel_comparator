magic
tech sky130A
timestamp 1621153998
<< checkpaint >>
rect -1853 -1878 2114 2081
<< error_p >>
rect 113 114 148 115
<< nwell >>
rect -261 100 799 810
<< mvnmos >>
rect -136 -114 -86 -14
rect 33 -114 83 -14
rect 257 -100 307 -50
rect 445 -214 495 -14
rect 549 -214 599 -14
rect 662 -214 712 -14
rect 131 -311 181 -261
rect -9 -429 91 -379
rect 131 -429 181 -379
rect 305 -568 355 -368
rect 445 -568 495 -368
<< mvpmos >>
rect -152 135 -52 235
rect -6 135 94 235
rect 257 135 307 735
rect 445 135 495 535
rect 549 135 599 535
rect 662 135 712 535
<< mvndiff >>
rect -208 -22 -136 -14
rect -208 -106 -191 -22
rect -162 -106 -136 -22
rect -208 -114 -136 -106
rect -86 -22 33 -14
rect -86 -106 -71 -22
rect 17 -106 33 -22
rect -86 -114 33 -106
rect 83 -22 153 -14
rect 83 -106 102 -22
rect 145 -106 153 -22
rect 405 -22 445 -14
rect 198 -100 257 -50
rect 307 -58 349 -50
rect 307 -92 323 -58
rect 341 -92 349 -58
rect 307 -100 349 -92
rect 83 -114 153 -106
rect 405 -206 413 -22
rect 431 -206 445 -22
rect 405 -214 445 -206
rect 495 -214 549 -14
rect 599 -22 662 -14
rect 599 -206 616 -22
rect 644 -206 662 -22
rect 599 -214 662 -206
rect 712 -22 756 -14
rect 712 -206 727 -22
rect 748 -206 756 -22
rect 712 -214 756 -206
rect 97 -269 131 -261
rect 97 -303 102 -269
rect 119 -303 131 -269
rect 97 -311 131 -303
rect 181 -272 234 -261
rect 181 -301 202 -272
rect 228 -301 234 -272
rect 181 -311 234 -301
rect 258 -376 305 -368
rect -57 -388 -9 -379
rect -57 -420 -48 -388
rect -26 -420 -9 -388
rect -57 -429 -9 -420
rect 91 -429 131 -379
rect 181 -387 221 -379
rect 181 -421 194 -387
rect 213 -421 221 -387
rect 181 -429 221 -421
rect 258 -557 269 -376
rect 295 -557 305 -376
rect 258 -568 305 -557
rect 355 -376 445 -368
rect 355 -560 372 -376
rect 430 -560 445 -376
rect 355 -568 445 -560
rect 495 -376 538 -368
rect 495 -560 510 -376
rect 530 -560 538 -376
rect 495 -568 538 -560
<< mvpdiff >>
rect -206 228 -152 235
rect -206 143 -194 228
rect -176 143 -152 228
rect -206 135 -152 143
rect -52 227 -6 235
rect -52 144 -43 227
rect -15 144 -6 227
rect -52 135 -6 144
rect 94 227 153 235
rect 94 143 117 227
rect 145 143 153 227
rect 94 135 153 143
rect 198 135 257 735
rect 307 725 433 735
rect 307 145 324 725
rect 422 535 433 725
rect 422 145 445 535
rect 307 135 445 145
rect 495 527 549 535
rect 495 143 512 527
rect 533 143 549 527
rect 495 135 549 143
rect 599 527 662 535
rect 599 142 612 527
rect 648 142 662 527
rect 599 135 662 142
rect 712 135 756 535
<< mvndiffc >>
rect -191 -106 -162 -22
rect -71 -106 17 -22
rect 102 -106 145 -22
rect 323 -92 341 -58
rect 413 -206 431 -22
rect 616 -206 644 -22
rect 727 -206 748 -22
rect 102 -303 119 -269
rect 202 -301 228 -272
rect -48 -420 -26 -388
rect 194 -421 213 -387
rect 269 -557 295 -376
rect 372 -560 430 -376
rect 510 -560 530 -376
<< mvpdiffc >>
rect -194 143 -176 228
rect -43 144 -15 227
rect 117 143 145 227
rect 324 145 422 725
rect 512 143 533 527
rect 612 142 648 527
<< mvpsubdiff >>
rect -232 -590 26 -576
rect -232 -697 -219 -590
rect 10 -697 26 -590
rect -232 -705 26 -697
<< mvnsubdiff >>
rect 464 770 760 776
rect 464 648 498 770
rect 733 648 760 770
rect 464 623 760 648
<< mvpsubdiffcont >>
rect -219 -697 10 -590
<< mvnsubdiffcont >>
rect 498 648 733 770
<< poly >>
rect 257 735 307 750
rect -152 235 -52 262
rect -6 235 94 262
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 445 535 495 558
rect 549 535 599 566
rect 662 535 712 558
rect -152 110 -52 135
rect -152 93 -144 110
rect -59 93 -52 110
rect -152 85 -52 93
rect -6 110 94 135
rect -6 93 2 110
rect 87 93 94 110
rect -6 85 94 93
rect 257 117 307 135
rect 296 86 307 117
rect 445 110 495 135
rect 445 49 453 110
rect 487 49 495 110
rect -136 -14 -86 -1
rect 33 -14 83 -1
rect 257 -50 307 27
rect 445 -14 495 49
rect 549 -14 599 135
rect 662 106 712 135
rect 662 12 670 106
rect 704 12 712 106
rect 662 -14 712 12
rect 257 -113 307 -100
rect -136 -201 -86 -114
rect 33 -132 83 -114
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect -136 -239 -86 -231
rect 131 -222 181 -215
rect 131 -239 139 -222
rect 173 -239 181 -222
rect 445 -227 495 -214
rect 549 -227 599 -214
rect 662 -228 712 -214
rect 131 -261 181 -239
rect 445 -303 495 -295
rect -9 -379 91 -355
rect 131 -379 181 -311
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 305 -368 355 -344
rect 445 -368 495 -343
rect -9 -454 91 -429
rect -9 -483 -1 -454
rect 71 -483 91 -454
rect 131 -462 181 -429
rect -9 -491 91 -483
rect 305 -593 355 -568
rect 445 -583 495 -568
rect 305 -618 313 -593
rect 347 -618 355 -593
rect 305 -627 355 -618
<< polycont >>
rect 557 566 591 596
rect -144 93 -59 110
rect 2 93 87 110
rect 257 86 296 117
rect 453 49 487 110
rect 670 12 704 106
rect 41 -170 71 -140
rect -128 -231 -94 -201
rect 139 -239 173 -222
rect 453 -343 487 -303
rect -1 -483 71 -454
rect 313 -618 347 -593
<< locali >>
rect -261 770 799 810
rect -261 758 498 770
rect -202 228 -167 235
rect -202 143 -194 228
rect -176 143 -167 228
rect -202 135 -167 143
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 109 227 153 235
rect 109 143 117 227
rect 145 143 153 227
rect 109 135 153 143
rect 198 135 249 735
rect 314 725 433 735
rect 314 145 324 725
rect 422 145 433 725
rect 464 648 498 758
rect 733 758 799 770
rect 733 648 760 758
rect 464 623 760 648
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 145
rect 504 527 541 535
rect 504 143 512 527
rect 533 143 541 527
rect 504 135 541 143
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 719 527 756 535
rect 719 143 727 527
rect 748 143 756 527
rect 719 135 756 143
rect -152 110 94 118
rect -152 93 -144 110
rect -59 93 2 110
rect 87 93 94 110
rect -152 85 94 93
rect 445 110 495 118
rect 445 49 453 110
rect 487 49 495 110
rect 445 41 495 49
rect 662 106 712 114
rect 662 12 670 106
rect 704 12 712 106
rect 662 4 712 12
rect -203 -22 -148 -14
rect -203 -106 -191 -22
rect -162 -106 -148 -22
rect -203 -114 -148 -106
rect -79 -22 25 -14
rect -79 -106 -71 -22
rect 17 -106 25 -22
rect -79 -114 25 -106
rect 94 -22 153 -14
rect 94 -106 102 -22
rect 145 -106 153 -22
rect 405 -22 439 -14
rect 315 -58 349 -50
rect 315 -92 323 -58
rect 341 -92 349 -58
rect 315 -100 349 -92
rect 94 -114 153 -106
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -201 -86 -193
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect 405 -206 413 -22
rect 431 -206 439 -22
rect 405 -214 439 -206
rect 608 -22 652 -14
rect 608 -206 616 -22
rect 644 -206 652 -22
rect 608 -214 652 -206
rect 719 -22 756 -14
rect 719 -206 727 -22
rect 748 -206 756 -22
rect 719 -214 756 -206
rect -136 -239 -86 -231
rect 131 -222 221 -215
rect 131 -239 139 -222
rect 173 -239 221 -222
rect 131 -244 221 -239
rect 185 -261 221 -244
rect 97 -269 125 -261
rect 97 -303 102 -269
rect 119 -303 125 -269
rect 97 -311 125 -303
rect 185 -272 234 -261
rect 185 -301 202 -272
rect 228 -301 234 -272
rect 185 -311 234 -301
rect 445 -303 495 -295
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect 258 -376 305 -368
rect -57 -388 -17 -379
rect -57 -420 -48 -388
rect -26 -420 -17 -388
rect -57 -429 -17 -420
rect 186 -387 221 -379
rect 186 -421 194 -387
rect 213 -421 221 -387
rect 186 -429 221 -421
rect -9 -454 79 -446
rect -9 -483 -1 -454
rect 71 -483 79 -454
rect -9 -491 79 -483
rect 258 -557 269 -376
rect 295 -557 305 -376
rect 258 -568 305 -557
rect 363 -376 438 -368
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
rect 503 -376 538 -368
rect 503 -560 510 -376
rect 530 -560 538 -376
rect 503 -568 538 -560
rect -232 -590 26 -576
rect -232 -697 -219 -590
rect 10 -647 26 -590
rect 305 -593 355 -585
rect 305 -618 313 -593
rect 347 -618 355 -593
rect 305 -627 355 -618
rect 10 -659 767 -647
rect 10 -697 25 -659
rect 53 -697 88 -659
rect 116 -697 153 -659
rect 181 -697 210 -659
rect 238 -697 273 -659
rect 301 -697 339 -659
rect 367 -697 396 -659
rect 424 -697 459 -659
rect 487 -697 518 -659
rect 546 -697 575 -659
rect 603 -697 638 -659
rect 666 -697 700 -659
rect 728 -697 767 -659
rect -232 -705 767 -697
<< viali >>
rect -194 143 -176 228
rect -43 144 -15 227
rect 117 143 145 227
rect 324 145 422 725
rect 557 566 591 596
rect 512 143 533 527
rect 612 142 648 527
rect 727 143 748 527
rect -144 93 -59 110
rect 2 93 87 110
rect 257 86 296 117
rect 453 49 487 110
rect 670 12 704 106
rect -191 -106 -162 -22
rect -71 -106 17 -22
rect 102 -106 145 -22
rect 323 -92 341 -58
rect 41 -170 71 -140
rect -128 -231 -94 -201
rect 413 -206 431 -22
rect 616 -206 644 -22
rect 727 -206 748 -22
rect 102 -303 119 -269
rect 202 -301 228 -272
rect 453 -343 487 -303
rect -48 -420 -26 -388
rect 194 -421 213 -387
rect -1 -483 71 -454
rect 269 -557 295 -376
rect 372 -560 430 -376
rect 510 -560 530 -376
rect 313 -618 347 -593
rect -219 -697 -191 -659
rect -162 -697 -134 -659
rect -99 -697 -71 -659
rect -32 -697 -4 -659
rect 25 -697 53 -659
rect 88 -697 116 -659
rect 153 -697 181 -659
rect 210 -697 238 -659
rect 273 -697 301 -659
rect 339 -697 367 -659
rect 396 -697 424 -659
rect 459 -697 487 -659
rect 518 -697 546 -659
rect 575 -697 603 -659
rect 638 -697 666 -659
rect 700 -697 728 -659
<< metal1 >>
rect -261 758 799 810
rect -203 228 -167 235
rect -203 143 -194 228
rect -176 143 -167 228
rect -203 118 -167 143
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 109 227 153 235
rect 109 143 117 227
rect 145 143 153 227
rect -203 110 94 118
rect -203 93 -144 110
rect -59 93 2 110
rect 87 93 94 110
rect -203 85 94 93
rect 109 117 153 143
rect -203 -22 -148 85
rect 109 -14 153 86
rect -203 -106 -191 -22
rect -162 -106 -148 -22
rect -203 -114 -148 -106
rect -79 -22 25 -14
rect -79 -106 -71 -22
rect 17 -106 25 -22
rect -79 -114 25 -106
rect 94 -22 153 -14
rect 94 -106 102 -22
rect 145 -106 153 -22
rect 94 -114 153 -106
rect 198 135 249 735
rect 314 725 433 735
rect 314 145 324 725
rect 422 145 433 725
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 145
rect 504 527 541 535
rect 504 143 512 527
rect 533 143 541 527
rect 504 135 541 143
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 719 527 756 535
rect 719 143 727 527
rect 748 143 756 527
rect 719 135 756 143
rect 198 72 243 135
rect -203 -528 -151 -114
rect -136 -201 -86 -193
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect -136 -239 -86 -231
rect -57 -388 -15 -114
rect 198 -125 243 41
rect 314 27 346 135
rect 257 -20 346 27
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 315 -58 349 -50
rect 315 -92 323 -58
rect 341 -92 349 -58
rect 33 -178 80 -170
rect 315 -182 349 -92
rect -57 -420 -48 -388
rect -26 -420 -15 -388
rect -57 -429 -15 -420
rect 97 -211 349 -182
rect 97 -269 126 -211
rect 363 -263 388 86
rect 445 110 495 118
rect 445 49 453 110
rect 487 49 495 110
rect 445 41 495 49
rect 509 114 541 135
rect 509 106 712 114
rect 509 14 670 106
rect 405 12 670 14
rect 704 12 712 106
rect 405 4 712 12
rect 405 -14 541 4
rect 727 -14 756 135
rect 405 -22 439 -14
rect 405 -206 413 -22
rect 431 -206 439 -22
rect 405 -228 439 -206
rect 608 -22 652 -14
rect 608 -206 616 -22
rect 644 -206 652 -22
rect 405 -249 591 -228
rect 97 -303 102 -269
rect 119 -303 126 -269
rect -9 -454 79 -446
rect -9 -483 -1 -454
rect 71 -483 79 -454
rect -9 -491 79 -483
rect 97 -647 126 -303
rect 196 -272 234 -266
rect 196 -301 202 -272
rect 228 -301 234 -272
rect 363 -279 538 -263
rect 196 -307 234 -301
rect 445 -303 495 -295
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect 509 -368 538 -279
rect 258 -376 305 -368
rect 186 -387 221 -379
rect 186 -421 194 -387
rect 220 -421 221 -387
rect 186 -429 221 -421
rect 258 -557 269 -376
rect 295 -557 305 -376
rect 258 -568 305 -557
rect 363 -376 438 -368
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
rect 503 -376 538 -368
rect 503 -560 510 -376
rect 530 -560 538 -376
rect 503 -568 538 -560
rect 561 -585 591 -249
rect 305 -593 591 -585
rect 305 -618 313 -593
rect 347 -618 591 -593
rect 305 -627 591 -618
rect 608 -647 652 -206
rect 719 -22 756 -14
rect 719 -206 727 -22
rect 748 -206 756 -22
rect 719 -214 756 -206
rect -232 -659 767 -647
rect -232 -697 -219 -659
rect -191 -697 -162 -659
rect -134 -697 -99 -659
rect -71 -697 -32 -659
rect -4 -697 25 -659
rect 53 -697 88 -659
rect 116 -697 153 -659
rect 181 -697 210 -659
rect 238 -697 273 -659
rect 301 -697 339 -659
rect 367 -697 396 -659
rect 424 -697 459 -659
rect 487 -697 518 -659
rect 546 -697 575 -659
rect 603 -697 638 -659
rect 666 -697 700 -659
rect 728 -697 767 -659
rect -232 -705 767 -697
<< via1 >>
rect -43 144 -15 227
rect 109 86 153 117
rect 324 145 422 725
rect 557 566 591 596
rect 612 142 648 527
rect 257 86 296 117
rect 198 41 243 72
rect -128 -231 -94 -201
rect 363 86 388 117
rect 41 -170 71 -140
rect 198 -165 243 -125
rect 453 49 487 110
rect -1 -483 71 -454
rect -203 -568 -151 -528
rect 202 -301 228 -272
rect 453 -343 487 -303
rect 194 -421 213 -387
rect 213 -421 220 -387
rect 221 -568 258 -528
rect 372 -560 430 -376
<< metal2 >>
rect -261 758 799 810
rect 314 725 433 735
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 314 145 324 725
rect 422 145 433 725
rect 549 603 846 648
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 145
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 153 86 257 117
rect 296 86 363 117
rect 445 110 495 118
rect 445 72 453 110
rect 243 49 453 72
rect 487 49 495 110
rect 243 41 495 49
rect -275 -140 80 -117
rect -275 -163 41 -140
rect 33 -170 41 -163
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -201 -86 -193
rect -136 -207 -128 -201
rect -361 -231 -128 -207
rect -94 -231 -86 -201
rect -361 -273 -86 -231
rect 246 -236 796 -235
rect 241 -261 796 -236
rect 196 -272 796 -261
rect 196 -301 202 -272
rect 228 -281 796 -272
rect 228 -301 266 -281
rect 196 -307 266 -301
rect 445 -303 495 -295
rect 196 -311 234 -307
rect 280 -327 431 -319
rect 221 -343 431 -327
rect 221 -355 300 -343
rect 221 -379 250 -355
rect 186 -387 250 -379
rect 186 -421 194 -387
rect 220 -421 250 -387
rect 186 -429 250 -421
rect 363 -368 431 -343
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect 363 -376 438 -368
rect -9 -454 79 -446
rect -9 -483 -1 -454
rect 71 -483 79 -454
rect -9 -491 79 -483
rect -151 -568 221 -528
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
<< via2 >>
rect -43 144 -15 227
rect 324 145 422 725
rect 612 142 648 527
rect 198 -165 243 -125
rect 453 -343 487 -303
rect -1 -483 71 -454
<< metal3 >>
rect -261 758 799 810
rect -261 -446 -226 758
rect -48 227 -10 758
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 314 725 433 758
rect 314 145 324 725
rect 422 145 433 725
rect 314 135 433 145
rect 604 527 656 758
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 243 -165 378 -125
rect 338 -295 378 -165
rect 338 -303 495 -295
rect 338 -338 453 -303
rect 445 -343 453 -338
rect 487 -343 495 -303
rect 445 -351 495 -343
rect -261 -454 79 -446
rect -261 -483 -1 -454
rect 71 -483 79 -454
rect -261 -491 79 -483
<< labels >>
rlabel viali 159 -678 159 -678 1 GND
rlabel metal2 816 632 816 632 1 EN
rlabel metal2 759 -262 759 -262 1 Ihyst
rlabel metal2 -340 -224 -340 -224 1 INN
rlabel metal2 -271 -159 -271 -159 1 INP
rlabel metal1 742 59 742 59 1 VOUT
<< end >>
