magic
tech sky130A
timestamp 1623667149
<< mvpsubdiff >>
rect 875 0 1075 25
<< locali >>
rect 875 0 1075 25
<< metal1 >>
rect 875 456 885 554
rect 1065 456 1075 554
rect -10 62 8 429
rect 875 176 1075 215
rect 1391 62 1435 429
rect 875 0 1075 25
<< via1 >>
rect 157 182 192 209
rect 332 182 367 209
<< metal2 >>
rect 151 209 198 215
rect 151 182 157 209
rect 192 182 198 209
rect 151 -12 198 182
rect 326 209 373 215
rect 326 182 332 209
rect 367 182 373 209
rect 326 -12 373 182
use inverter3v3  inverter3v3_3
timestamp 1623667149
transform 1 0 525 0 1 0
box 0 0 175 554
use inverter3v3  inverter3v3_2
timestamp 1623667149
transform 1 0 350 0 1 0
box 0 0 175 554
use inverter3v3  inverter3v3_1
timestamp 1623667149
transform 1 0 175 0 1 0
box 0 0 175 554
use inverter3v3  inverter3v3_0
timestamp 1623667149
transform 1 0 0 0 1 0
box 0 0 175 554
use inverter3v3  inverter3v3_4
timestamp 1623667149
transform 1 0 700 0 1 0
box 0 0 175 554
use inverter3v3  inverter3v3_5
timestamp 1623667149
transform 1 0 1075 0 1 0
box 0 0 175 554
use inverter3v3  inverter3v3_6
timestamp 1623667149
transform 1 0 1250 0 1 0
box 0 0 175 554
<< labels >>
rlabel metal1 1433 187 1433 187 7 OUT
rlabel metal1 969 8 969 8 1 GND
rlabel metal1 1069 492 1069 492 1 VCC
rlabel metal1 881 487 881 487 1 VADJ
rlabel metal2 178 -7 178 -7 1 OUT1
rlabel metal2 348 -5 348 -5 1 OUT2
rlabel metal1 -7 186 -7 186 3 IN
<< end >>
