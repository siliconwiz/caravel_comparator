magic
tech sky130A
timestamp 1621157240
<< nwell >>
rect -261 102 799 810
rect -261 100 243 102
rect 445 100 799 102
<< mvnmos >>
rect -136 -114 -86 -14
rect 33 -114 83 -14
rect 257 -100 307 -50
rect 445 -214 495 -14
rect 549 -214 599 -14
rect 662 -214 712 -14
rect 131 -311 181 -261
rect -9 -429 91 -379
rect 131 -429 181 -379
rect 305 -568 355 -368
rect 445 -568 495 -368
<< mvpmos >>
rect -152 135 -52 235
rect -6 135 94 235
rect 257 135 307 735
rect 445 135 495 535
rect 549 135 599 535
rect 662 135 712 535
<< mvndiff >>
rect -208 -22 -136 -14
rect -208 -106 -191 -22
rect -162 -106 -136 -22
rect -208 -114 -136 -106
rect -86 -22 33 -14
rect -86 -106 -71 -22
rect 17 -106 33 -22
rect -86 -114 33 -106
rect 83 -22 153 -14
rect 83 -106 102 -22
rect 145 -106 153 -22
rect 405 -22 445 -14
rect 198 -58 257 -50
rect 198 -92 206 -58
rect 235 -92 257 -58
rect 198 -100 257 -92
rect 307 -58 349 -50
rect 307 -92 323 -58
rect 341 -92 349 -58
rect 307 -100 349 -92
rect 83 -114 153 -106
rect 405 -206 413 -22
rect 431 -206 445 -22
rect 405 -214 445 -206
rect 495 -214 549 -14
rect 599 -22 662 -14
rect 599 -206 616 -22
rect 644 -206 662 -22
rect 599 -214 662 -206
rect 712 -22 756 -14
rect 712 -206 727 -22
rect 748 -206 756 -22
rect 712 -214 756 -206
rect 97 -269 131 -261
rect 97 -303 102 -269
rect 119 -303 131 -269
rect 97 -311 131 -303
rect 181 -272 234 -261
rect 181 -301 202 -272
rect 228 -301 234 -272
rect 181 -311 234 -301
rect 258 -376 305 -368
rect -57 -388 -9 -379
rect -57 -420 -48 -388
rect -26 -420 -9 -388
rect -57 -429 -9 -420
rect 91 -387 131 -379
rect 91 -421 102 -387
rect 119 -421 131 -387
rect 91 -429 131 -421
rect 181 -387 221 -379
rect 181 -421 194 -387
rect 213 -421 221 -387
rect 181 -429 221 -421
rect 258 -557 269 -376
rect 295 -557 305 -376
rect 258 -568 305 -557
rect 355 -376 445 -368
rect 355 -560 372 -376
rect 430 -560 445 -376
rect 355 -568 445 -560
rect 495 -376 538 -368
rect 495 -560 510 -376
rect 530 -560 538 -376
rect 495 -568 538 -560
<< mvpdiff >>
rect 204 727 257 735
rect -206 228 -152 235
rect -206 143 -194 228
rect -176 143 -152 228
rect -206 135 -152 143
rect -52 227 -6 235
rect -52 144 -43 227
rect -15 144 -6 227
rect -52 135 -6 144
rect 94 227 153 235
rect 94 143 117 227
rect 145 143 153 227
rect 94 135 153 143
rect 204 143 212 727
rect 241 143 257 727
rect 204 135 257 143
rect 307 727 433 735
rect 307 143 322 727
rect 425 535 433 727
rect 425 143 445 535
rect 307 135 445 143
rect 495 527 549 535
rect 495 143 512 527
rect 532 143 549 527
rect 495 135 549 143
rect 599 527 662 535
rect 599 142 612 527
rect 648 142 662 527
rect 599 135 662 142
rect 712 527 756 535
rect 712 143 727 527
rect 748 143 756 527
rect 712 135 756 143
<< mvndiffc >>
rect -191 -106 -162 -22
rect -71 -106 17 -22
rect 102 -106 145 -22
rect 206 -92 235 -58
rect 323 -92 341 -58
rect 413 -206 431 -22
rect 616 -206 644 -22
rect 727 -206 748 -22
rect 102 -303 119 -269
rect 202 -301 228 -272
rect -48 -420 -26 -388
rect 102 -421 119 -387
rect 194 -421 213 -387
rect 269 -557 295 -376
rect 372 -560 430 -376
rect 510 -560 530 -376
<< mvpdiffc >>
rect -194 143 -176 228
rect -43 144 -15 227
rect 117 143 145 227
rect 212 143 241 727
rect 322 143 425 727
rect 512 143 532 527
rect 612 142 648 527
rect 727 143 748 527
<< mvpsubdiff >>
rect 575 -308 767 -294
rect -232 -522 221 -511
rect -232 -697 -219 -522
rect 208 -647 221 -522
rect 575 -647 587 -308
rect 208 -659 587 -647
rect 208 -697 238 -659
rect 546 -697 587 -659
rect 755 -697 767 -308
rect -232 -705 767 -697
<< mvnsubdiff >>
rect -228 751 143 768
rect -228 357 -205 751
rect 123 357 143 751
rect 499 761 742 768
rect -228 337 143 357
rect 499 685 535 761
rect 728 685 742 761
rect 499 665 742 685
<< mvpsubdiffcont >>
rect -219 -697 208 -522
rect 238 -697 546 -659
rect 587 -697 755 -308
<< mvnsubdiffcont >>
rect -205 357 123 751
rect 535 685 728 761
<< poly >>
rect 257 735 307 750
rect -152 235 -52 262
rect -6 235 94 262
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 445 535 495 558
rect 549 535 599 566
rect 662 535 712 558
rect -152 110 -52 135
rect -152 93 -144 110
rect -59 93 -52 110
rect -152 85 -52 93
rect -6 110 94 135
rect -6 93 2 110
rect 87 93 94 110
rect -6 85 94 93
rect 257 110 307 135
rect 257 88 265 110
rect 299 88 307 110
rect 257 80 307 88
rect 445 110 495 135
rect 445 49 453 110
rect 487 49 495 110
rect 257 19 307 27
rect -136 -14 -86 -1
rect 33 -14 83 -1
rect 257 -12 266 19
rect 299 -12 307 19
rect 257 -50 307 -12
rect 445 -14 495 49
rect 549 -14 599 135
rect 662 106 712 135
rect 662 12 670 106
rect 704 12 712 106
rect 662 -14 712 12
rect 257 -113 307 -100
rect -136 -201 -86 -114
rect 33 -132 83 -114
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect -136 -239 -86 -231
rect 131 -222 181 -215
rect 131 -239 139 -222
rect 173 -239 181 -222
rect 445 -227 495 -214
rect 549 -227 599 -214
rect 662 -228 712 -214
rect 131 -261 181 -239
rect 445 -303 495 -295
rect -9 -379 91 -355
rect 131 -379 181 -311
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 305 -368 355 -344
rect 445 -368 495 -343
rect -9 -454 91 -429
rect -9 -483 -1 -454
rect 71 -483 91 -454
rect 131 -462 181 -429
rect -9 -491 91 -483
rect 305 -593 355 -568
rect 445 -583 495 -568
rect 305 -618 313 -593
rect 347 -618 355 -593
rect 305 -627 355 -618
<< polycont >>
rect 557 566 591 596
rect -144 93 -59 110
rect 2 93 87 110
rect 265 88 299 110
rect 453 49 487 110
rect 266 -12 299 19
rect 670 12 704 106
rect 41 -170 71 -140
rect -128 -231 -94 -201
rect 139 -239 173 -222
rect 453 -343 487 -303
rect -1 -483 71 -454
rect 313 -618 347 -593
<< locali >>
rect -261 799 799 810
rect -261 769 198 799
rect 756 769 799 799
rect -261 761 799 769
rect -261 758 535 761
rect -261 751 170 758
rect -261 357 -205 751
rect 123 357 170 751
rect -261 309 170 357
rect 50 308 170 309
rect 204 727 249 735
rect -202 228 -167 235
rect -202 143 -194 228
rect -176 143 -167 228
rect -202 135 -167 143
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 109 227 153 235
rect 109 143 117 227
rect 145 143 153 227
rect 109 135 153 143
rect 204 143 212 727
rect 241 143 249 727
rect 204 135 249 143
rect 314 727 433 735
rect 314 143 322 727
rect 425 143 433 727
rect 468 685 535 758
rect 728 685 799 761
rect 468 631 799 685
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 143
rect 504 527 540 535
rect 504 143 512 527
rect 532 143 540 527
rect 504 135 540 143
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 719 527 756 535
rect 719 143 727 527
rect 748 143 756 527
rect 719 135 756 143
rect -152 110 94 118
rect -152 93 -144 110
rect -59 93 2 110
rect 87 93 94 110
rect -152 85 94 93
rect 257 110 307 118
rect 257 88 265 110
rect 299 88 307 110
rect 257 80 307 88
rect 445 110 495 118
rect 445 49 453 110
rect 487 49 495 110
rect 445 41 495 49
rect 662 106 712 114
rect 257 19 307 27
rect 257 -12 266 19
rect 299 -12 307 19
rect 662 12 670 106
rect 704 12 712 106
rect 662 4 712 12
rect -203 -22 -148 -14
rect -203 -106 -191 -22
rect -162 -106 -148 -22
rect -203 -114 -148 -106
rect -79 -22 25 -14
rect -79 -106 -71 -22
rect 17 -106 25 -22
rect -79 -114 25 -106
rect 94 -22 153 -14
rect 257 -20 307 -12
rect 94 -106 102 -22
rect 145 -106 153 -22
rect 405 -22 439 -14
rect 198 -58 243 -50
rect 198 -92 206 -58
rect 235 -92 243 -58
rect 198 -100 243 -92
rect 315 -58 349 -50
rect 315 -92 323 -58
rect 341 -92 349 -58
rect 315 -100 349 -92
rect 94 -114 153 -106
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -201 -86 -193
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect 405 -206 413 -22
rect 431 -206 439 -22
rect 405 -214 439 -206
rect 608 -22 652 -14
rect 608 -206 616 -22
rect 644 -206 652 -22
rect 608 -214 652 -206
rect 719 -22 756 -14
rect 719 -206 727 -22
rect 748 -206 756 -22
rect 719 -214 756 -206
rect -136 -239 -86 -231
rect 131 -222 221 -215
rect 131 -239 139 -222
rect 173 -239 221 -222
rect 131 -244 221 -239
rect 185 -261 221 -244
rect 97 -269 125 -261
rect 97 -303 102 -269
rect 119 -303 125 -269
rect 97 -311 125 -303
rect 185 -272 234 -261
rect 185 -301 202 -272
rect 228 -301 234 -272
rect 185 -311 234 -301
rect 445 -303 495 -295
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect 575 -308 767 -294
rect 258 -376 305 -368
rect -57 -388 -17 -379
rect -57 -420 -48 -388
rect -26 -420 -17 -388
rect -57 -429 -17 -420
rect 97 -387 126 -379
rect 97 -421 102 -387
rect 119 -421 126 -387
rect -9 -454 79 -446
rect -9 -483 -1 -454
rect 71 -483 79 -454
rect -9 -491 79 -483
rect 97 -511 126 -421
rect 186 -387 221 -379
rect 186 -421 194 -387
rect 213 -421 221 -387
rect 186 -429 221 -421
rect -232 -522 221 -511
rect -232 -697 -219 -522
rect 208 -647 221 -522
rect 258 -557 269 -376
rect 295 -557 305 -376
rect 258 -568 305 -557
rect 363 -376 438 -368
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
rect 503 -376 538 -368
rect 503 -560 510 -376
rect 530 -560 538 -376
rect 503 -568 538 -560
rect 305 -593 355 -585
rect 305 -618 313 -593
rect 347 -618 355 -593
rect 305 -627 355 -618
rect 575 -647 587 -308
rect 208 -659 587 -647
rect 208 -697 210 -659
rect 546 -697 575 -659
rect 755 -697 767 -308
rect -232 -705 767 -697
<< viali >>
rect 198 769 756 799
rect -204 358 123 751
rect -194 143 -176 228
rect -43 144 -15 227
rect 117 143 145 227
rect 212 143 241 727
rect 322 143 425 727
rect 557 566 591 596
rect 512 143 532 527
rect 612 142 648 527
rect 727 143 748 527
rect -144 93 -59 110
rect 2 93 87 110
rect 265 88 299 110
rect 453 49 487 110
rect 266 -12 299 19
rect 670 12 704 106
rect -191 -106 -162 -22
rect -71 -106 17 -22
rect 102 -106 145 -22
rect 206 -92 235 -58
rect 323 -92 341 -58
rect 41 -170 71 -140
rect -128 -231 -94 -201
rect 413 -206 431 -22
rect 616 -206 644 -22
rect 727 -206 748 -22
rect 102 -303 119 -269
rect 202 -301 228 -272
rect 453 -343 487 -303
rect -48 -420 -26 -388
rect 102 -421 119 -387
rect -1 -483 71 -454
rect 194 -421 213 -387
rect 269 -557 295 -376
rect 372 -560 430 -376
rect 510 -560 530 -376
rect 313 -618 347 -593
rect -219 -697 -191 -659
rect -162 -697 -134 -659
rect -99 -697 -71 -659
rect -32 -697 -4 -659
rect 25 -697 53 -659
rect 88 -697 116 -659
rect 153 -697 181 -659
rect 210 -697 238 -659
rect 273 -697 301 -659
rect 339 -697 367 -659
rect 396 -697 424 -659
rect 459 -697 487 -659
rect 518 -697 546 -659
rect 575 -697 587 -659
rect 587 -697 603 -659
rect 638 -697 666 -659
rect 700 -697 728 -659
<< metal1 >>
rect -261 799 799 810
rect -261 769 198 799
rect 756 769 799 799
rect -261 758 799 769
rect -261 751 170 758
rect -261 358 -204 751
rect 123 358 170 751
rect -261 309 170 358
rect 50 308 170 309
rect 204 727 249 735
rect -203 228 -167 235
rect -203 143 -194 228
rect -176 143 -167 228
rect -203 118 -167 143
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 109 227 153 235
rect 109 143 117 227
rect 145 143 153 227
rect -203 110 94 118
rect -203 93 -144 110
rect -59 93 2 110
rect 87 93 94 110
rect -203 85 94 93
rect 109 117 153 143
rect 204 143 212 727
rect 241 143 249 727
rect 204 135 249 143
rect 314 727 433 735
rect 314 143 322 727
rect 425 143 433 727
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 143
rect 504 527 541 535
rect 504 143 512 527
rect 532 143 541 527
rect 504 135 541 143
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 719 527 756 535
rect 719 143 727 527
rect 748 143 756 527
rect 719 135 756 143
rect 109 110 388 117
rect 109 88 265 110
rect 299 88 388 110
rect -203 -22 -148 85
rect 109 80 388 88
rect 109 -14 153 80
rect -203 -106 -191 -22
rect -162 -106 -148 -22
rect -203 -114 -148 -106
rect -79 -22 25 -14
rect -79 -106 -71 -22
rect 17 -106 25 -22
rect -79 -114 25 -106
rect 94 -22 153 -14
rect 263 19 307 27
rect 263 -12 266 19
rect 299 -12 307 19
rect 263 -20 307 -12
rect 94 -106 102 -22
rect 145 -106 153 -22
rect 198 -58 243 -50
rect 198 -92 206 -58
rect 235 -92 243 -58
rect 198 -100 243 -92
rect 315 -58 349 -50
rect 315 -92 323 -58
rect 341 -92 349 -58
rect 94 -114 153 -106
rect -203 -528 -151 -114
rect -57 -163 -15 -114
rect 33 -140 80 -132
rect 33 -170 41 -140
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -201 -86 -193
rect -136 -231 -128 -201
rect -94 -231 -86 -201
rect -136 -239 -86 -231
rect -57 -388 -15 -178
rect 315 -182 349 -92
rect -57 -420 -48 -388
rect -26 -420 -15 -388
rect -57 -429 -15 -420
rect 97 -211 349 -182
rect 97 -269 126 -211
rect 363 -263 388 80
rect 445 110 495 118
rect 445 49 453 110
rect 487 49 495 110
rect 445 41 495 49
rect 509 114 541 135
rect 509 106 712 114
rect 509 14 670 106
rect 405 12 670 14
rect 704 12 712 106
rect 405 4 712 12
rect 405 -14 541 4
rect 727 -14 756 135
rect 405 -22 439 -14
rect 405 -206 413 -22
rect 431 -206 439 -22
rect 405 -228 439 -206
rect 608 -22 652 -14
rect 608 -206 616 -22
rect 644 -206 652 -22
rect 405 -249 591 -228
rect 97 -303 102 -269
rect 119 -303 126 -269
rect 97 -387 126 -303
rect 196 -272 234 -266
rect 196 -301 202 -272
rect 228 -301 234 -272
rect 363 -279 538 -263
rect 196 -307 234 -301
rect 445 -303 495 -295
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect 509 -368 538 -279
rect 258 -376 305 -368
rect 97 -421 102 -387
rect 119 -421 126 -387
rect 97 -429 126 -421
rect 186 -387 221 -379
rect 186 -421 194 -387
rect 220 -421 221 -387
rect 186 -429 221 -421
rect -9 -454 79 -446
rect -9 -483 -1 -454
rect 71 -483 79 -454
rect -9 -491 79 -483
rect 258 -528 269 -376
rect -203 -557 269 -528
rect 295 -557 305 -376
rect -203 -568 305 -557
rect 363 -376 438 -368
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
rect 503 -376 538 -368
rect 503 -560 510 -376
rect 530 -560 538 -376
rect 503 -568 538 -560
rect 561 -585 591 -249
rect 305 -593 591 -585
rect 305 -618 313 -593
rect 347 -618 591 -593
rect 305 -627 591 -618
rect 608 -294 652 -206
rect 719 -22 756 -14
rect 719 -206 727 -22
rect 748 -206 756 -22
rect 719 -214 756 -206
rect 608 -647 767 -294
rect -232 -659 767 -647
rect -232 -697 -219 -659
rect -191 -697 -162 -659
rect -134 -697 -99 -659
rect -71 -697 -32 -659
rect -4 -697 25 -659
rect 53 -697 88 -659
rect 116 -697 153 -659
rect 181 -697 210 -659
rect 238 -697 273 -659
rect 301 -697 339 -659
rect 367 -697 396 -659
rect 424 -697 459 -659
rect 487 -697 518 -659
rect 546 -697 575 -659
rect 603 -697 638 -659
rect 666 -697 700 -659
rect 728 -697 767 -659
rect -232 -705 767 -697
<< via1 >>
rect 198 769 756 799
rect -204 358 123 751
rect -43 144 -15 227
rect 212 143 241 727
rect 322 143 425 727
rect 557 566 591 596
rect 612 142 648 527
rect 266 -12 299 19
rect 206 -92 235 -58
rect 41 -170 71 -140
rect -128 -231 -94 -201
rect 453 49 487 110
rect 202 -301 228 -272
rect 453 -343 487 -303
rect 194 -421 213 -387
rect 213 -421 220 -387
rect -1 -483 71 -454
rect 372 -560 430 -376
<< metal2 >>
rect -261 799 799 810
rect -261 769 198 799
rect 756 769 799 799
rect -261 758 799 769
rect -261 751 170 758
rect -261 358 -204 751
rect 123 358 170 751
rect -261 309 170 358
rect 50 308 170 309
rect 204 727 249 735
rect -48 227 -10 235
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 204 143 212 727
rect 241 143 249 727
rect 204 135 249 143
rect 314 727 433 735
rect 314 143 322 727
rect 425 143 433 727
rect 549 603 846 648
rect 549 596 599 603
rect 549 566 557 596
rect 591 566 599 596
rect 549 558 599 566
rect 314 135 433 143
rect 604 527 656 535
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect -361 -122 -226 85
rect 204 72 243 135
rect 445 110 495 118
rect 445 72 453 110
rect 204 49 453 72
rect 487 49 495 110
rect 204 41 495 49
rect 204 -50 243 41
rect 257 19 307 27
rect 257 -12 266 19
rect 299 -12 307 19
rect 257 -20 307 -12
rect 198 -58 243 -50
rect 198 -92 206 -58
rect 235 -92 243 -58
rect 198 -100 243 -92
rect -361 -140 80 -122
rect -361 -163 41 -140
rect 33 -170 41 -163
rect 71 -170 80 -140
rect 33 -178 80 -170
rect -136 -201 -86 -193
rect -136 -208 -128 -201
rect -361 -231 -128 -208
rect -94 -231 -86 -201
rect -361 -277 -86 -231
rect 246 -236 796 -235
rect 241 -261 796 -236
rect 196 -272 796 -261
rect -361 -462 -226 -277
rect 196 -301 202 -272
rect 228 -281 796 -272
rect 228 -301 266 -281
rect 196 -307 266 -301
rect 445 -303 495 -295
rect 196 -311 234 -307
rect 280 -327 431 -319
rect 221 -343 431 -327
rect 221 -355 300 -343
rect 221 -379 250 -355
rect 186 -387 250 -379
rect 186 -421 194 -387
rect 220 -421 250 -387
rect 186 -429 250 -421
rect 363 -368 431 -343
rect 445 -343 453 -303
rect 487 -343 495 -303
rect 445 -351 495 -343
rect 363 -376 438 -368
rect -9 -454 79 -446
rect -9 -483 -1 -454
rect 71 -483 79 -454
rect -9 -491 79 -483
rect 363 -560 372 -376
rect 430 -560 438 -376
rect 363 -568 438 -560
<< via2 >>
rect 198 769 756 799
rect -204 358 123 751
rect -43 144 -15 227
rect 322 143 425 727
rect 612 142 648 527
rect 266 -12 299 19
rect 206 -92 235 -58
rect 453 -343 487 -303
rect -1 -483 71 -454
<< metal3 >>
rect -261 799 799 810
rect -261 769 198 799
rect 756 769 799 799
rect -261 758 799 769
rect -261 751 170 758
rect -261 358 -204 751
rect 123 358 170 751
rect -261 309 170 358
rect -261 -446 -226 309
rect -48 227 -10 309
rect 50 308 170 309
rect 314 727 433 758
rect -48 144 -43 227
rect -15 144 -10 227
rect -48 135 -10 144
rect 314 143 322 727
rect 425 143 433 727
rect 314 135 433 143
rect 604 527 656 758
rect 604 142 612 527
rect 648 142 656 527
rect 604 135 656 142
rect 314 27 353 135
rect 257 19 353 27
rect 257 -12 266 19
rect 299 -12 353 19
rect 257 -20 353 -12
rect 198 -58 243 -50
rect 198 -92 206 -58
rect 235 -92 243 -58
rect 198 -125 243 -92
rect 198 -165 378 -125
rect 338 -295 378 -165
rect 338 -303 495 -295
rect 338 -338 453 -303
rect 445 -343 453 -338
rect 487 -343 495 -303
rect 445 -351 495 -343
rect -261 -454 79 -446
rect -261 -483 -1 -454
rect 71 -483 79 -454
rect -261 -491 79 -483
<< labels >>
rlabel viali 159 -678 159 -678 1 GND
rlabel metal2 816 632 816 632 1 EN
rlabel metal2 759 -262 759 -262 1 Ihyst
rlabel metal2 -340 -224 -340 -224 1 INN
rlabel metal2 -271 -159 -271 -159 1 INP
rlabel metal1 742 59 742 59 1 VOUT
<< end >>
